//------------------------------------------------------------------------
//    final_top.sv Spring 2020                                          --
//    Adapted from lab8.sv, lab8                                        --
//    Toplevel                                                          --
//------------------------------------------------------------------------


module final_top 
(   
    input               CLOCK_50,
    input        [3:0]  KEY,         //bit 0 is set up as Reset
    output logic [6:0]  HEX0, HEX1,
    //// VGA Interface ////
    output logic [7:0]  VGA_R, VGA_G, VGA_B, //VGA RGB
    output logic VGA_CLK,           //VGA Clock
                    VGA_SYNC_N,        //VGA Sync signal
                    VGA_BLANK_N,       //VGA Blank signal
                    VGA_VS,            //VGA virtical sync signal
                    VGA_HS,            //VGA horizontal sync signal
    //// CY7C67200 Interface ////
    inout  wire  [15:0] OTG_DATA,   //CY7C67200 Data bus 16 Bits
    output logic [1:0]  OTG_ADDR,   //CY7C67200 Address 2 Bits
    output logic        OTG_CS_N,   //CY7C67200 Chip Select
                        OTG_RD_N,   //CY7C67200 Write
                        OTG_WR_N,   //CY7C67200 Read
                        OTG_RST_N,  //CY7C67200 Reset
    input               OTG_INT,    //CY7C67200 Interrupt
    //// SDRAM Interface for Nios II Software ////
    output logic [12:0] DRAM_ADDR,  //SDRAM Address 13 Bits
    inout  wire  [31:0] DRAM_DQ,    //SDRAM Data 32 Bits
    output logic [1:0]  DRAM_BA,    //SDRAM Bank Address 2 Bits
    output logic [3:0]  DRAM_DQM,   //SDRAM Data Mast 4 Bits
    output logic        DRAM_RAS_N, //SDRAM Row Address Strobe
                        DRAM_CAS_N, //SDRAM Column Address Strobe
                        DRAM_CKE,   //SDRAM Clock Enable
                        DRAM_WE_N,  //SDRAM Write Enable
                        DRAM_CS_N,  //SDRAM Chip Select
                        DRAM_CLK,   //SDRAM Clock
    //// WM8731 Audio Interface ////
    input        [17:0] SW, 
    output logic [17:0] LEDR,
    inout  wire         I2C_SDAT,
    output logic        I2C_SCLK, AUD_XCK, AUD_BCLK, AUD_DACLRCK, AUD_DACDAT
);
    
    logic Reset_h, Clk;
    logic [7:0] keycode;
    logic [9:0] DrawX, DrawY;
    logic [11:0] frame_counter;
    logic [9:0] GroundY, StickmanTop;
    logic is_stickman, is_ground, is_coin, is_score, is_star, is_human, is_win_text, is_lose_text, is_select_text;
    
    logic coin_collide;
    logic [4:0] status;  // {selecting, waiting, playing, win, lose}
    logic [1:0] level_status; // 01 = level 1; 10 = level 2
    logic restart;
    assign restart = status[3];


    logic [9:0] CoinY[3];
    logic [12:0] CoinFrameX[3];
    logic [2:0] CoinStatus;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    

    //////// Interface between NIOS II and EZ-OTG chip ////////
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
    
    hpi_io_intf hpi_io_inst(
        .Clk(Clk), .Reset(Reset_h),
        // signals connected to NIOS II
        .from_sw_address(hpi_addr), .from_sw_data_in(hpi_data_in), .from_sw_data_out(hpi_data_out),
        .from_sw_r(hpi_r), .from_sw_w(hpi_w), .from_sw_cs(hpi_cs), .from_sw_reset(hpi_reset),
        // signals connected to EZ-OTG chip
        .OTG_DATA(OTG_DATA), .OTG_ADDR(OTG_ADDR), .OTG_RD_N(OTG_RD_N),    
        .OTG_WR_N(OTG_WR_N), .OTG_CS_N(OTG_CS_N), .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     lab8_soc m_lab8_soc(
        .clk_clk(Clk), .reset_reset_n(1'b1),    // Never reset NIOS
        .sdram_wire_addr(DRAM_ADDR), .sdram_wire_ba(DRAM_BA), .sdram_wire_cas_n(DRAM_CAS_N),
        .sdram_wire_cke(DRAM_CKE), .sdram_wire_cs_n(DRAM_CS_N), .sdram_wire_dq(DRAM_DQ),   
        .sdram_wire_dqm(DRAM_DQM), .sdram_wire_ras_n(DRAM_RAS_N), .sdram_wire_we_n(DRAM_WE_N), .sdram_c1k_clk(DRAM_CLK),
        .keycode_export(keycode),  
        .otg_hpi_address_export(hpi_addr), .otg_hpi_data_in_port(hpi_data_in), .otg_hpi_data_out_port(hpi_data_out),
        .otg_hpi_cs_export(hpi_cs), .otg_hpi_r_export(hpi_r), .otg_hpi_w_export(hpi_w), .otg_hpi_reset_export(hpi_reset)
    );
    

    //////// VGA control and interface ////////

    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    
    VGA_controller vga_controller_instance(
        .*,                 // Clk, VGA_HS, VGA_VS, VGA_BLANK_N, VGA_SYNC_N
        .Reset(Reset_h), .VGA_CLK, .DrawX, .DrawY	// Active-high reset, 25 MHz VGA clock input, XY coordinates
	);
    // Which signal should be frame_clk? --> "One way to keep track of frames is simply by keeping track of tile Vertical Sync (vs) signal"


    stickman my_stickman (
        .*,                 // Clk, DrawX, DrawY, is_stickman, keycode, GroundY, playing
        .Reset(Reset_h), .frame_clk(VGA_VS) // Active-high reset, The clock indicating a new frame (~60Hz)
	);

    background  my_background ( 
        .*,                 // Clk, DrawX, DrawY, is_ground, is_coin, keycode, CoinFrameX[3], CoinY[3], CoinStatus, GroundY, playing, frame_counter
        .Reset(Reset_h), .frame_clk(VGA_VS)	// Active-high reset, The clock indicating a new frame (~60Hz)
    );

    score       my_score(.*, .Reset(Reset_h));  // Clk, DrawX, DrawY, is_score, is_board, frame_counter, Active-high reset
    star        my_star (.*, .Reset(Reset_h));  // Clk, DrawX, DrawY, CoinStatus, is_star, frame_counter, Active-high reset
    
    human       my_human (.*, .Reset(Reset_h)); // Clk ,DrawX,DrawY, is_human, Active-high reset
    win_text    my_win   (.*, .Reset(Reset_h)); // Clk, DrawX, DrawY, is_win_text, Active-high reset
    lose_text   my_lose  (.*, .Reset(Reset_h)); // Clk, DrawX, DrawY, is_lose_text, Active-high reset
    select_text my_select(.*, .Reset(Reset_h)); // Clk, DrawX, DrawY, is_lose_text, Active-high reset

    color_mapper color_instance(.*); 	// is_stickman, is_ground, is_coin, is_coin, is_board, DrawX, DrawY, VGA_R, VGA_G, VGA_B, status

    game_logic logic_instance(  
        .*,                     // Clk, keycode, status, StickmanBottom, GroundY, CoinFrameX[3], CoinY[3], CoinStatus, frame_counter
        .Reset(Reset_h), .frame_clk(VGA_VS)     // Active-high reset, The clock indicating a new frame (~60Hz)
    );

    
    // Display keycode on hex display
    HexDriver hex_inst_0 (keycode[3:0], HEX0);
    HexDriver hex_inst_1 (keycode[7:4], HEX1);


    ///////// Audio Control ////////
    Sound_Top Sound_Top_inst( 
        .clk(Clk), .reset(KEY[0]), .SoundSelect({coin_collide, status[1:0]}),
        .SDIN(I2C_SDAT), .SCLK(I2C_SCLK), .USB_clk(AUD_XCK), .BCLK(AUD_BCLK),
        .DAC_LR_CLK(AUD_DACLRCK), .DAC_DATA(AUD_DACDAT), .ACK_LEDR(LEDR[2:0])
    );
    
endmodule